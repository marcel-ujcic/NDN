library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VAJA2_1 is
    Port ( pick : in STD_LOGIC_VECTOR(1 downto 0);
			  a : in  STD_LOGIC;
           b : in  STD_LOGIC;
			  c : in  STD_LOGIC;
			  d : in  STD_LOGIC;
           f : out  STD_LOGIC);
end VAJA2_1;

architecture Behavioral of VAJA2_1 is
	 
begin
	
	


end Behavioral;

