----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:41:56 04/28/2021 
-- Design Name: 
-- Module Name:    mux2_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2_1 is
    Port ( in_0,in_1 : in  STD_LOGIC_VECTOR (1 downto 0);
           mux_select : in  STD_LOGIC;
           mux_out : out  STD_LOGIC_VECTOR (1 downto 0));
end mux2_1;

architecture Behavioral of mux2_1 is

begin
	
	mux_out <= in_0 when mux_select = '0' else in_1; 


end Behavioral;

